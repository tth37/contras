@Head
NAME Not
INPUT a
OUTPUT out
SYMBOL NAND NAND1
@Body
NAND1(a = a, b = a) => (out = na)
@End
OUTPUT out = na

import And from "And.cdl"

@Head
NAME And4
INPUT a[3:0]
OUTPUT out
SYMBOL And And1, And2, And3

@Body
And1(a = a[0], b = a[1]) => (out = a01)
And2(a = a[2], b = a[3]) => (out = a23)
And3(a = a01, b = a23) => (out = res)

@End
OUTPUT out = res

# .\contras.exe .\And4.cdl .\test\And4.in .\test\And4.out
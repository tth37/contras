import And4 from "And4.cdl"
import Not from "Not.cdl"

@Head
NAME DMux2Way4
INPUT a, b, D
OUTPUT Y3, Y2, Y1, Y0
SYMBOL And4 And41, And42, And43, And44
SYMBOL Not Not1, Not2

@Body
Not1(a=a)=>(out=na)
Not2(a=b)=>(out=nb)
And41(a[0]=D, a[1]=D, a[2]=na, a[3]=nb)=>(out=W0)
And42(a[0]=D, a[1]=D, a[2]=a, a[3]=nb)=>(out=W1)
And43(a[0]=D, a[1]=D, a[2]=na, a[3]=b)=>(out=W2)
And44(a[0]=D, a[1]=D, a[2]=a, a[3]=b)=>(out=W3)

@End
OUTPUT Y0=W0,Y1=W1, Y2=W2, Y3=W3
@Head
NAME RSFlipFlop
INPUT R, S
OUTPUT Q, NQ
STATE SQ = 0, SNQ = 1
SYMBOL NAND NAND1, NAND2
@Body
NAND1(a = S, b = SNQ) => (out = t1)
NAND2(a = R, b = SQ) => (out = t2)
@End
STATE SQ = t1, SNQ = t2
OUTPUT Q = t1, NQ = t2

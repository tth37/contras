@Head
NAME Not
INPUT a
OUTPUT out
SYMBOL NAND Nand1

@Body
Nand1(a = a, b = a) => (out = res)

@End
OUTPUT out = res

# .\contras.exe .\Not.cdl .\test\Not.in .\test\Not.out
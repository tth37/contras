import And4 from "And4.cdl"
import Not from "Not.cdl"
import And from "And.cdl"

@Head
NAME Mux4Way1
INPUT a, b
INPUT D0, D1, D2, D3
OUTPUT W, NW
SYMBOL And And1, And2, And3, And4
SYMBOL And4 And41
SYMBOL NAND NAND1, NAND2, NAND3, NAND4
SYMBOL Not Not1, Not2, Not3

@Body
Not1(a=a)=>(out=na)
Not2(a=b)=>(out=nb)
And1(a=na, b=nb)=>(out=nanb)
And2(a=a, b=nb)=>(out=anb)
And3(a=na, b=b)=>(out=nab)
And4(a=a, b=b)=>(out=ab)
NAND1(a=nanb, b=D0)=>(out=d0)
NAND2(a=anb, b=D1)=>(out=d1)
NAND3(a=nab, b=D2)=>(out=d2)
NAND4(a=ab, b=D3)=>(out=d3)
And41(a[0]=d0, a[1]=d1, a[2]=d2, a[3]=d3)=>(out=nresult)
Not3(a=nresult)=>(out=result)

@End
OUTPUT W=result, NW=nresult

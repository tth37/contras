import Not from "Not.cdl"
@Head
NAME And
INPUT a, b
OUTPUT out
SYMBOL NAND NAND1
SYMBOL Not Not1
@Body
NAND1(a = a, b = b) => (out = nab)
Not1(a = nab) => (out = ab)
@End
OUTPUT out = ab

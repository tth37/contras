import And4 from "And4.cdl"
import Not from "Not.cdl"
import And from "And.cdl"

@Head
NAME Mux8Way1
INPUT c, b, a
INPUT D0, D1, D2, D3, D4, D5, D6, D7
OUTPUT W, NW
SYMBOL And And1
SYMBOL And4 And41, And42, And43, And44, And45, And46, And47, And48, And49, And410
SYMBOL Not Not1, Not2, Not3, Not4, Not5, Not6, Not7, Not8, Not9, Not10, Not11, Not12

@Body
Not1(a=a)=>(out=na)
Not2(a=b)=>(out=nb)
Not3(a=c)=>(out=nc)
And41(a[0]=nc, a[1]=nb, a[2]=na, a[3]=D0)=>(out=d0)
And42(a[0]=nc, a[1]=nb, a[2]=a, a[3]=D1)=>(out=d1)
And43(a[0]=nc, a[1]=b, a[2]=na, a[3]=D2)=>(out=d2)
And44(a[0]=nc, a[1]=b, a[2]=a, a[3]=D3)=>(out=d3)
And45(a[0]=c, a[1]=nb, a[2]=na, a[3]=D4)=>(out=d4)
And46(a[0]=c, a[1]=nb, a[2]=a, a[3]=D5)=>(out=d5)
And47(a[0]=c, a[1]=b, a[2]=na, a[3]=D6)=>(out=d6)
And48(a[0]=c, a[1]=b, a[2]=a, a[3]=D7)=>(out=d7)
Not5(a=d0)=>(out=nD0)
Not6(a=d1)=>(out=nD1)
Not7(a=d2)=>(out=nD2)
Not8(a=d3)=>(out=nD3)
Not9(a=d4)=>(out=nD4)
Not10(a=d5)=>(out=nD5)
Not11(a=d6)=>(out=nD6)
Not12(a=d7)=>(out=nD7)
And49(a[0]=nD0, a[1]=nD1, a[2]=nD2, a[3]=nD3)=>(out=nD0123)
And410(a[0]=nD4, a[1]=nD5, a[2]=nD6, a[3]=nD7)=>(out=nD4567)
And1(a=nD0123, b=nD4567)=>(out=nresult)
Not4(a=nresult)=>(out=result)

@End
OUTPUT W=result, NW=nresult